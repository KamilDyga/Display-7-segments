library ieee;

use ieee.std_logic_1164.all;

entity decoder is
	port(
		
		digit		: in std_logic_vector(3 downto 0);
		segment	: out std_logic_vector(6 downto 0)
	
	);
end decoder;
	
architecture basic of decoder is

begin
	
	--std_logic_vector(to_unsigned(10, 8))
	--segment(6 downto 0) <= 	"1111110" when digit = "0000" else
	--								"0110000" when digit = "0001" else
	--								"1101101" when digit = "0010" else
	--								"1111001" when digit = "0011" else
	--								"0110011" when digit = "0100" else
	--								"1011011" when digit = "0101" else
	--								"1011111" when digit = "0110" else
	--								"0000001";
									-- uzupełnić inne cyfry, napisać testbench
	with digit select
		segment (6 downto 0) <=	 "1111110" when "0000", --0
										 "0110000" when "0001", --1
										 "1101101" when "0010", --2
										 "1111001" when "0011", --3
										 "0110011" when "0100", --4
										 "1011011" when "0101", --5
										 "1011111" when "0110", --6
										 "1110000" when "0111", --7
										 "1111111" when "1000", --8
										 "1111011" when "1001", --9
										 "1110111" when "1010", --A
										 "0011111" when "1011", --B
										 "1001110" when "1100", --C
										 "0111101" when "1101", --D
										 "1001111" when "1110", --E
										 "1000111" when "1111", --F
										 "0000001" when others ;
			
end basic;